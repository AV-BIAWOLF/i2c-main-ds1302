// params.vh

`ifndef params
`define params

    parameter WRITE_TEST_COUNT = 2;
    parameter READ_TEST_COUNT = 2;
    parameter CLK_PERIOD = 10;

`endif